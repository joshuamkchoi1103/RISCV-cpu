// Code your testbench here
// or browse Examples
//`include "run.do"
//`include "milestone2_quicktest_tb.sv"
//`include "test.sv"
//`include "fix2flt_tb.sv"
//`include "flt2fix_tb.sv"
`include "fltflt_no_rnd_tb.sv"